module sva (
   spi_slave_inter.dut Spi_slave_test_vif
);
    endmodule